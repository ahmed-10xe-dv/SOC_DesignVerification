// Interface to connect to DUT
interface AndGateInterface();
  logic [3:0] input_a, input_b;
  logic [3:0] output_res;  
endinterface