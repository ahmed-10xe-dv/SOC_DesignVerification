// Interface to connect to DUT
interface CounterInterface();
  logic  clk,rst, up, load ;
  logic [7:0] loadin, y;  
endinterface