
// Interface to connect to DUT
interface AndGateInterface();
    logic A, B, C, D;   // Inputs for the 4-input AND gate
    logic Y;            // Output result  
  endinterface